library verilog;
use verilog.vl_types.all;
entity ramtest is
end ramtest;

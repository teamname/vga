library verilog;
use verilog.vl_types.all;
entity r_tb is
end r_tb;

library verilog;
use verilog.vl_types.all;
entity vga_driver_tb is
end vga_driver_tb;

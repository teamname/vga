library verilog;
use verilog.vl_types.all;
entity Rom is
end Rom;

library verilog;
use verilog.vl_types.all;
entity duck_hunt_tb is
end duck_hunt_tb;
